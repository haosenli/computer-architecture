/*
 * EE469 Autumn 2022
 * Haosen Li, Peter Tran
 * 
 * This file computes or-ing bits together.
 *
 * Inputs:
 * A - 1 bit, A bit.
 * B - 1 bit, B bit.
 * sel - 1 bit, selects the out value.
 *
 * Outputs:
 * Cout - 1 bit, Output of A or B.
 */
module orAB (
	input logic A, B, sel,
	output logic out
	);
	
	logic or1;
	
	// A or B
	or #5 or_AB (or1, A, B);
	
	// Mux to decide whether to output A or B or 0
	mux_2x1 mux2x1 (.in({or1, 1'b0}), .sel(sel), .out(out)); 
	
endmodule