module data_id(
	input 
	);

	
endmodule
