/*
 * EE469 Autumn 2022
 * Haosen Li, Peter Tran
 * 
 * This file contains the adder controller file.
 *
 * Inputs:
 * ctrl - 3 bits, Control signal.
 *
 * Outputs:
 * 
 */

module adder_controller(
        input  logic [2:0] ctrl
    );